`timescale 1 ns / 1 ps

module stream_slave_test (
   output logic M_AXIS_TREADY
);
   
   initial M_AXIS_TREADY = 1;

endmodule 
